/* Роутер содержит в себе внутренний буфер, с количеством ячеек, равному
 * количеству процессоров (CPU_N), и размером равном размеру сообщения
 * (MSG_SIZE).
 * Каждый процессор (с номером id) может оставить сообщение, переданное по своему
 * выделенному каналу (data[id]) для процессора, номер которого передан также по 
 * выделенному каналу (addr[id]), установив свою линию записи (we[id]).
 * Аналогичным образом каждый процессор может считать по своей линии данные
 * для процессора с адресом addr.
 */

module sm_router
(
	input clk,
	inout [MSG_SIZE-1:0] data[CPU_N-1:0], /* линия данных - по 1 на каждый процессор */
	input addr[CPU_N-1:0], /* линия выбора адреса для чтения / записи по 1 на каждый проц */
	input we[CPU_N-1:0], /* линия бита записи по 1 на каждый проц. если нет сигнала, значит чтение */
	input [3:0] id /* id процессора, который обращается к роутеру */
);
	parameter CPU_N = 4;
	parameter MSG_SIZE = 32;
	reg [MSG_SIZE-1:0] internal_data[CPU_N-1];

	always @(posedge clk)
	begin
		if (we[id])
			internal_data[addr] <= data[id];
		else	
			data[id] <= internal_data[addr];
	end
endmodule
